library ieee;
use ieee.std_logic_1164.all;

entity i2c_controller_tb_rd is
end entity i2c_controller_tb_rd;

architecture sim of i2c_controller_tb_rd is
  constant TB_SYSTEM_CLK_FREQUENCY : integer := 20e6;
  constant TB_SYSTEM_CLK_PERIOD : time := 1000 ms / TB_SYSTEM_CLK_FREQUENCY;
  constant TB_I2C_BUS_KBITPS : integer := 100000;
  signal tb_sda : std_logic := 'H';
  signal tb_scl : std_logic := 'H';
  signal tb_clk : std_logic := '0';
  signal tb_nena : std_logic := '0';
  signal tb_rw : std_logic := '1';
  signal tb_data_out : std_logic_vector(7 downto 0);
  signal tb_data_in : std_logic_vector(7 downto 0) := x"51";
  signal tb_address : std_logic_vector(6 downto 0) := "1001001";
begin

  UUT: entity work.i2c_controller(rtl)
  generic map (
    SYSTEM_CLK_FREQUENCY => TB_SYSTEM_CLK_FREQUENCY,
    I2C_BUS_KBITPS => TB_I2C_BUS_KBITPS
  )
  port map (
    sda => to_x01(tb_sda),
    scl => to_x01(tb_scl),
    clk => tb_clk,
    nena => tb_nena,
    rw => tb_rw,
    data_out => tb_data_out,
    data_in => tb_data_in,
    address => tb_address
  );

  tb_clk <= not tb_clk after TB_SYSTEM_CLK_PERIOD / 2;
  tb_sda <= 'H';
  tb_scl <= 'H';
  
  process
  begin
    wait for 195000 ns;
    tb_nena <= '1';
    wait;
  end process;
  
  ack: process
  begin
    wait for 89925 ns;
    tb_sda <= '0';
    wait for 10000 ns;
    tb_sda <= 'H';
    wait;
  end process;

end architecture sim;